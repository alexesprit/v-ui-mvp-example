module main

import gui

fn main() {
	v := gui.create_app_view()
	v.start()
}
