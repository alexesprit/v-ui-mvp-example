module main

import view

fn main() {
	v := view.create_view()
	v.run()
}
