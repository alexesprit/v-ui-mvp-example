module view

pub interface IAppView {
	set_textbox_value(value int)
}
